--
-- VHDL Architecture ece411.IR3regsplitter.untitled
--
-- Created:
--          by - adalton2.ews (gelib-057-40.ews.illinois.edu)
--          at - 23:16:50 04/16/14
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY IR3regsplitter IS
-- Declarations

END IR3regsplitter ;

--
ARCHITECTURE untitled OF IR3regsplitter IS
BEGIN
END ARCHITECTURE untitled;

